library verilog;
use verilog.vl_types.all;
entity CombinedASU2_vlg_check_tst is
    port(
        leds1           : in     vl_logic;
        leds2           : in     vl_logic;
        leds3           : in     vl_logic;
        leds4           : in     vl_logic;
        leds5           : in     vl_logic;
        leds6           : in     vl_logic;
        leds7           : in     vl_logic;
        leds21          : in     vl_logic;
        leds22          : in     vl_logic;
        leds23          : in     vl_logic;
        leds24          : in     vl_logic;
        leds25          : in     vl_logic;
        leds26          : in     vl_logic;
        leds27          : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end CombinedASU2_vlg_check_tst;
